`timescale 1ns / 1ps


module pbg_tb;

reg a,b,c,d;

wire e;

pbg u_test(
.a(a ),
.b(b ),
.c(c ),
.d(d ),

.e(e )
);

initial begin
    a = 1'b0;
    b = 1'b0;
    c = 1'b0;
    d = 1'b0;
end

always@(a or b or c or d) begin
    a <= #60 ~a;
    b <= #100 ~b;
    c <= #150 ~c;
    d <= #200 ~d;
end

initial begin
    #1000
    $finish;
end



endmodule